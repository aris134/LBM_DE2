library verilog;
use verilog.vl_types.all;
entity tb_display is
end tb_display;
