module tb_display;
	initial begin
		$display("Testing....");
	end
endmodule
