module LBM_DE2	#(GRID_DIM=16,
		DATA_WIDTH=32)(
		
		input CLOCK_50,
		input RESET);

endmodule
